module ex62_top(  
KEY,  
CLOCK_50,  
HEX0,HEX1,HEX2,HEX3,HEX4  
);  
   
//INPUT AND OUTPUT declare independently  
  input [1:0] KEY;  
  input CLOCK_50;  
  output [6:0] HEX0;  
  output [6:0]HEX1;  
  output [6:0]HEX2;  
  output [6:0]HEX3;  
  output [6:0]HEX4;  
   
  wire [15:0] count;   
  wire [3:0] BCD0,BCD1,BCD2,BCD3,BCD4;  
  wire tick;  
  wire en;  
  
  clkdiv_50000 ck0(CLOCK_50,tick); 
  assign en = ~KEY[0]&tick; 
   
  counter_16 B1(CLOCK_50,en,~KEY[1],count);  
  bin2bcd_16 B2(count,BCD0,BCD1,BCD2,BCD3,BCD4);  
   
  hex_to_7seg reg0(HEX0,BCD0);  
  hex_to_7seg reg1(HEX1,BCD1);  
  hex_to_7seg reg2(HEX2,BCD2);  
  hex_to_7seg reg3(HEX3,BCD3);  
  hex_to_7seg reg4(HEX4,BCD4);  
   
endmodule  