//------------------------------
// Module name: allpass processor
// Function: Simply to pass input to output
// Creator:  Peter Cheung
// Version:  1.1
// Date:     24 Jan 2014
//------------------------------

module processor (sysclk, data_in, data_out,data_valid);

   input          data_valid;
	input				sysclk;		// system clock
	input [9:0]		data_in;		// 10-bit input data
	output [9:0] 	data_out;	// 10-bit output data

	wire				sysclk;
	wire [9:0]		data_in;
	reg [9:0] 		data_out;
	wire [9:0]		x,y,z;
	wire           full,pulse;
	reg            q;

	parameter 		ADC_OFFSET = 10'h181; //385
	parameter 		DAC_OFFSET = 10'h200; //512

	assign x = data_in[9:0] - ADC_OFFSET;		// x is input in 2's complement
	
	pulse_gen p(pulse,data_valid,sysclk);
	FIFO fifo(sysclk,x[9:0],rdreq,pulse,full,z[9:0]);
	always @(posedge sysclk)
	    q <=full;
		 
	assign rdreq = q & data_valid;
	assign y =x[9:0]+{z[9],z[9:1]};
	 
	//  Now clock y output with system clock
	always @(posedge sysclk)
		data_out <=  y + DAC_OFFSET;
		
endmodule
	